module E300ArtyDevKit
(
    input  logic        cpu_ext_clk,
    input  logic        cpu_clock,
    input  logic        cpu_rst_n,

    input  logic        jtag_rst_n,
    input  logic        jtag_tck,
    input  logic        jtag_tms,
    input  logic        jtag_tdi,
    output logic        jtag_tdo,

    inout  logic [31:0] gpios,

    output logic        qspi_sck,
    output logic        qspi_cs,
    inout  logic [3:0]  qspi_dq
);

    logic [31:0]        gpio_oe, gpio_ival, gpio_oval;
    logic [3:0]         qspi_dq_oe, qspi_dq_ival, qspi_dq_oval;

    // Drive GPIO and SPI pins
    generate
    // GPIO
    for(genvar i = 0; i < 32; i++) begin
        assign gpios[i] = gpio_oe[i] ? gpio_oval[i] : 1'bZ;
    end
    assign gpio_ival = gpios;
    // QSPI
    for (genvar j = 0; j < 4; j++) begin
        assign qspi_dq[j] = qspi_dq_oe[j] ? qspi_dq_oval[j] : 1'bZ;
    end
    assign qspi_dq_ival = qspi_dq;
    endgenerate

    // Core
    E300ArtyDevKitPlatform E300ArtyDevKitPlatform_inst
    (
        .clock                            (cpu_clock        ),
        .reset                            (1'b0             ),

        .io_pins_aon_erst_n_i_ival        (cpu_rst_n        ),
        .io_pins_aon_erst_n_i_po          (/* UNCONNECTED */),
        .io_pins_aon_erst_n_o_oval        (/* UNCONNECTED */),
        .io_pins_aon_erst_n_o_oe          (/* UNCONNECTED */),
        .io_pins_aon_erst_n_o_ie          (/* UNCONNECTED */),
        .io_pins_aon_erst_n_o_poe         (/* UNCONNECTED */),
        .io_pins_aon_erst_n_o_pue         (/* UNCONNECTED */),
        .io_pins_aon_erst_n_o_ds          (/* UNCONNECTED */),
        .io_pins_aon_erst_n_o_ds1         (/* UNCONNECTED */),
        .io_pins_aon_erst_n_o_ps          (/* UNCONNECTED */),
        .io_pins_aon_lfextclk_i_ival      (cpu_ext_clk      ),
        .io_pins_aon_lfextclk_i_po        (/* UNCONNECTED */),
        .io_pins_aon_lfextclk_o_oval      (/* UNCONNECTED */),
        .io_pins_aon_lfextclk_o_oe        (/* UNCONNECTED */),
        .io_pins_aon_lfextclk_o_ie        (/* UNCONNECTED */),
        .io_pins_aon_lfextclk_o_pue       (/* UNCONNECTED */),
        .io_pins_aon_lfextclk_o_poe       (/* UNCONNECTED */),
        .io_pins_aon_lfextclk_o_ps        (/* UNCONNECTED */),
        .io_pins_aon_lfextclk_o_ds        (/* UNCONNECTED */),
        .io_pins_aon_lfextclk_o_ds1       (/* UNCONNECTED */),
        .io_pins_aon_pmu_dwakeup_n_i_ival (1'b0             ),
        .io_pins_aon_pmu_dwakeup_n_i_po   (/* UNCONNECTED */),
        .io_pins_aon_pmu_dwakeup_n_o_oval (/* UNCONNECTED */),
        .io_pins_aon_pmu_dwakeup_n_o_oe   (/* UNCONNECTED */),
        .io_pins_aon_pmu_dwakeup_n_o_ie   (/* UNCONNECTED */),
        .io_pins_aon_pmu_dwakeup_n_o_pue  (/* UNCONNECTED */),
        .io_pins_aon_pmu_dwakeup_n_o_ps   (/* UNCONNECTED */),
        .io_pins_aon_pmu_dwakeup_n_o_ds   (/* UNCONNECTED */),
        .io_pins_aon_pmu_dwakeup_n_o_ds1  (/* UNCONNECTED */),
        .io_pins_aon_pmu_vddpaden_i_ival  (1'b0             ),
        .io_pins_aon_pmu_vddpaden_i_po    (/* UNCONNECTED */),
        .io_pins_aon_pmu_vddpaden_o_oval  (/* UNCONNECTED */),
        .io_pins_aon_pmu_vddpaden_o_oe    (/* UNCONNECTED */),
        .io_pins_aon_pmu_vddpaden_o_ie    (/* UNCONNECTED */),
        .io_pins_aon_pmu_vddpaden_o_pue   (/* UNCONNECTED */),
        .io_pins_aon_pmu_dwakeup_n_o_poe  (/* UNCONNECTED */),
        .io_pins_aon_pmu_vddpaden_o_ps    (/* UNCONNECTED */),
        .io_pins_aon_pmu_vddpaden_o_ds    (/* UNCONNECTED */),
        .io_pins_aon_pmu_vddpaden_o_ds1   (/* UNCONNECTED */),
        .io_pins_aon_pmu_vddpaden_o_poe   (/* UNCONNECTED */),

        .io_jtag_reset                    (~jtag_rst_n      ),
        .io_pins_jtag_TCK_i_ival          (jtag_tck         ),
        .io_pins_jtag_TCK_i_po            (/* UNCONNECTED */),
        .io_pins_jtag_TCK_o_oval          (/* UNCONNECTED */),
        .io_pins_jtag_TCK_o_oe            (/* UNCONNECTED */),
        .io_pins_jtag_TCK_o_ie            (/* UNCONNECTED */),
        .io_pins_jtag_TMS_i_ival          (jtag_tms         ),
        .io_pins_jtag_TMS_i_po            (/* UNCONNECTED */),
        .io_pins_jtag_TMS_o_oval          (/* UNCONNECTED */),
        .io_pins_jtag_TMS_o_oe            (/* UNCONNECTED */),
        .io_pins_jtag_TMS_o_ie            (/* UNCONNECTED */),
        .io_pins_jtag_TDI_i_ival          (jtag_tdi         ),
        .io_pins_jtag_TDI_i_po            (/* UNCONNECTED */),
        .io_pins_jtag_TDI_o_oval          (/* UNCONNECTED */),
        .io_pins_jtag_TDI_o_oe            (/* UNCONNECTED */),
        .io_pins_jtag_TDI_o_ie            (/* UNCONNECTED */),
        .io_pins_jtag_TDO_i_ival          (1'b0             ),
        .io_pins_jtag_TDO_i_po            (/* UNCONNECTED */),
        .io_pins_jtag_TDO_o_oval          (jtag_tdo         ),
        .io_pins_jtag_TDO_o_oe            (/* UNCONNECTED */),
        .io_pins_jtag_TDO_o_ie            (/* UNCONNECTED */),

        .io_pins_gpio_pins_0_i_ival       (gpio_ival[0]     ),
        .io_pins_gpio_pins_0_i_po         (/* UNCONNECTED */),
        .io_pins_gpio_pins_0_o_oval       (gpio_oval[0]     ),
        .io_pins_gpio_pins_0_o_oe         (gpio_oe[0]       ),
        .io_pins_gpio_pins_0_o_ie         (/* UNCONNECTED */),
        .io_pins_gpio_pins_1_i_ival       (gpio_ival[1]     ),
        .io_pins_gpio_pins_1_i_po         (/* UNCONNECTED */),
        .io_pins_gpio_pins_1_o_oval       (gpio_oval[1]     ),
        .io_pins_gpio_pins_1_o_oe         (gpio_oe[1]       ),
        .io_pins_gpio_pins_1_o_ie         (/* UNCONNECTED */),
        .io_pins_gpio_pins_2_i_ival       (gpio_ival[2]     ),
        .io_pins_gpio_pins_2_i_po         (/* UNCONNECTED */),
        .io_pins_gpio_pins_2_o_oval       (gpio_oval[2]     ),
        .io_pins_gpio_pins_2_o_oe         (gpio_oe[2]       ),
        .io_pins_gpio_pins_2_o_ie         (/* UNCONNECTED */),
        .io_pins_gpio_pins_3_i_ival       (gpio_ival[3]     ),
        .io_pins_gpio_pins_3_i_po         (/* UNCONNECTED */),
        .io_pins_gpio_pins_3_o_oval       (gpio_oval[3]     ),
        .io_pins_gpio_pins_3_o_oe         (gpio_oe[3]       ),
        .io_pins_gpio_pins_3_o_ie         (/* UNCONNECTED */),
        .io_pins_gpio_pins_4_i_ival       (gpio_ival[4]     ),
        .io_pins_gpio_pins_4_i_po         (/* UNCONNECTED */),
        .io_pins_gpio_pins_4_o_oval       (gpio_oval[4]     ),
        .io_pins_gpio_pins_4_o_oe         (gpio_oe[4]       ),
        .io_pins_gpio_pins_4_o_ie         (/* UNCONNECTED */),
        .io_pins_gpio_pins_5_i_ival       (gpio_ival[5]     ),
        .io_pins_gpio_pins_5_i_po         (/* UNCONNECTED */),
        .io_pins_gpio_pins_5_o_oval       (gpio_oval[5]     ),
        .io_pins_gpio_pins_5_o_oe         (gpio_oe[5]       ),
        .io_pins_gpio_pins_5_o_ie         (/* UNCONNECTED */),
        .io_pins_gpio_pins_6_i_ival       (gpio_ival[6]     ),
        .io_pins_gpio_pins_6_i_po         (/* UNCONNECTED */),
        .io_pins_gpio_pins_6_o_oval       (gpio_oval[6]     ),
        .io_pins_gpio_pins_6_o_oe         (gpio_oe[6]       ),
        .io_pins_gpio_pins_6_o_ie         (/* UNCONNECTED */),
        .io_pins_gpio_pins_7_i_ival       (gpio_ival[7]     ),
        .io_pins_gpio_pins_7_i_po         (/* UNCONNECTED */),
        .io_pins_gpio_pins_7_o_oval       (gpio_oval[7]     ),
        .io_pins_gpio_pins_7_o_oe         (gpio_oe[7]       ),
        .io_pins_gpio_pins_7_o_ie         (/* UNCONNECTED */),
        .io_pins_gpio_pins_8_i_ival       (gpio_ival[8]     ),
        .io_pins_gpio_pins_8_i_po         (/* UNCONNECTED */),
        .io_pins_gpio_pins_8_o_oval       (gpio_oval[8]     ),
        .io_pins_gpio_pins_8_o_oe         (gpio_oe[8]       ),
        .io_pins_gpio_pins_8_o_ie         (/* UNCONNECTED */),
        .io_pins_gpio_pins_9_i_ival       (gpio_ival[9]     ),
        .io_pins_gpio_pins_9_i_po         (/* UNCONNECTED */),
        .io_pins_gpio_pins_9_o_oval       (gpio_oval[9]     ),
        .io_pins_gpio_pins_9_o_oe         (gpio_oe[9]       ),
        .io_pins_gpio_pins_9_o_ie         (/* UNCONNECTED */),
        .io_pins_gpio_pins_10_i_ival      (gpio_ival[10]    ),
        .io_pins_gpio_pins_10_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_10_o_oval      (gpio_oval[10]    ),
        .io_pins_gpio_pins_10_o_oe        (gpio_oe[10]      ),
        .io_pins_gpio_pins_10_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_11_i_ival      (gpio_ival[11]    ),
        .io_pins_gpio_pins_11_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_11_o_oval      (gpio_oval[11]    ),
        .io_pins_gpio_pins_11_o_oe        (gpio_oe[11]      ),
        .io_pins_gpio_pins_11_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_12_i_ival      (gpio_ival[12]    ),
        .io_pins_gpio_pins_12_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_12_o_oval      (gpio_oval[12]    ),
        .io_pins_gpio_pins_12_o_oe        (gpio_oe[12]      ),
        .io_pins_gpio_pins_12_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_13_i_ival      (gpio_ival[13]    ),
        .io_pins_gpio_pins_13_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_13_o_oval      (gpio_oval[13]    ),
        .io_pins_gpio_pins_13_o_oe        (gpio_oe[13]      ),
        .io_pins_gpio_pins_13_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_14_i_ival      (gpio_ival[14]    ),
        .io_pins_gpio_pins_14_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_14_o_oval      (gpio_oval[14]    ),
        .io_pins_gpio_pins_14_o_oe        (gpio_oe[14]      ),
        .io_pins_gpio_pins_14_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_15_i_ival      (gpio_ival[15]    ),
        .io_pins_gpio_pins_15_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_15_o_oval      (gpio_oval[15]    ),
        .io_pins_gpio_pins_15_o_oe        (gpio_oe[15]      ),
        .io_pins_gpio_pins_15_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_16_i_ival      (gpio_ival[16]    ),
        .io_pins_gpio_pins_16_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_16_o_oval      (gpio_oval[16]    ),
        .io_pins_gpio_pins_16_o_oe        (gpio_oe[16]      ),
        .io_pins_gpio_pins_16_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_17_i_ival      (gpio_ival[17]    ),
        .io_pins_gpio_pins_17_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_17_o_oval      (gpio_oval[17]    ),
        .io_pins_gpio_pins_17_o_oe        (gpio_oe[17]      ),
        .io_pins_gpio_pins_17_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_18_i_ival      (gpio_ival[18]    ),
        .io_pins_gpio_pins_18_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_18_o_oval      (gpio_oval[18]    ),
        .io_pins_gpio_pins_18_o_oe        (gpio_oe[18]      ),
        .io_pins_gpio_pins_18_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_19_i_ival      (gpio_ival[19]    ),
        .io_pins_gpio_pins_19_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_19_o_oval      (gpio_oval[19]    ),
        .io_pins_gpio_pins_19_o_oe        (gpio_oe[19]      ),
        .io_pins_gpio_pins_19_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_20_i_ival      (gpio_ival[20]    ),
        .io_pins_gpio_pins_20_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_20_o_oval      (gpio_oval[20]    ),
        .io_pins_gpio_pins_20_o_oe        (gpio_oe[20]      ),
        .io_pins_gpio_pins_20_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_21_i_ival      (gpio_ival[21]    ),
        .io_pins_gpio_pins_21_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_21_o_oval      (gpio_oval[21]    ),
        .io_pins_gpio_pins_21_o_oe        (gpio_oe[21]      ),
        .io_pins_gpio_pins_21_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_22_i_ival      (gpio_ival[22]    ),
        .io_pins_gpio_pins_22_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_22_o_oval      (gpio_oval[22]    ),
        .io_pins_gpio_pins_22_o_oe        (gpio_oe[22]      ),
        .io_pins_gpio_pins_22_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_23_i_ival      (gpio_ival[23]    ),
        .io_pins_gpio_pins_23_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_23_o_oval      (gpio_oval[23]    ),
        .io_pins_gpio_pins_23_o_oe        (gpio_oe[23]      ),
        .io_pins_gpio_pins_23_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_24_i_ival      (gpio_ival[24]    ),
        .io_pins_gpio_pins_24_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_24_o_oval      (gpio_oval[24]    ),
        .io_pins_gpio_pins_24_o_oe        (gpio_oe[24]      ),
        .io_pins_gpio_pins_24_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_25_i_ival      (gpio_ival[25]    ),
        .io_pins_gpio_pins_25_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_25_o_oval      (gpio_oval[25]    ),
        .io_pins_gpio_pins_25_o_oe        (gpio_oe[25]      ),
        .io_pins_gpio_pins_25_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_26_i_ival      (gpio_ival[26]    ),
        .io_pins_gpio_pins_26_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_26_o_oval      (gpio_oval[26]    ),
        .io_pins_gpio_pins_26_o_oe        (gpio_oe[26]      ),
        .io_pins_gpio_pins_26_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_27_i_ival      (gpio_ival[27]    ),
        .io_pins_gpio_pins_27_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_27_o_oval      (gpio_oval[27]    ),
        .io_pins_gpio_pins_27_o_oe        (gpio_oe[27]      ),
        .io_pins_gpio_pins_27_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_28_i_ival      (gpio_ival[28]    ),
        .io_pins_gpio_pins_28_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_28_o_oval      (gpio_oval[28]    ),
        .io_pins_gpio_pins_28_o_oe        (gpio_oe[28]      ),
        .io_pins_gpio_pins_28_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_29_i_ival      (gpio_ival[29]    ),
        .io_pins_gpio_pins_29_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_29_o_oval      (gpio_oval[29]    ),
        .io_pins_gpio_pins_29_o_oe        (gpio_oe[29]      ),
        .io_pins_gpio_pins_29_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_30_i_ival      (gpio_ival[30]    ),
        .io_pins_gpio_pins_30_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_30_o_oval      (gpio_oval[30]    ),
        .io_pins_gpio_pins_30_o_oe        (gpio_oe[30]      ),
        .io_pins_gpio_pins_30_o_ie        (/* UNCONNECTED */),
        .io_pins_gpio_pins_31_i_ival      (gpio_ival[31]    ),
        .io_pins_gpio_pins_31_i_po        (/* UNCONNECTED */),
        .io_pins_gpio_pins_31_o_oval      (gpio_oval[31]    ),
        .io_pins_gpio_pins_31_o_oe        (gpio_oe[31]      ),
        .io_pins_gpio_pins_31_o_ie        (/* UNCONNECTED */),

        .io_pins_qspi_sck_i_ival          (1'b0             ),
        .io_pins_qspi_sck_i_po            (/* UNCONNECTED */),
        .io_pins_qspi_sck_o_oval          (qspi_sck         ),
        .io_pins_qspi_sck_o_oe            (/* UNCONNECTED */),
        .io_pins_qspi_sck_o_ie            (/* UNCONNECTED */),
        .io_pins_qspi_cs_0_i_ival         (1'b0             ),
        .io_pins_qspi_cs_0_i_po           (/* UNCONNECTED */),
        .io_pins_qspi_cs_0_o_oval         (qspi_cs          ),
        .io_pins_qspi_cs_0_o_oe           (/* UNCONNECTED */),
        .io_pins_qspi_cs_0_o_ie           (/* UNCONNECTED */),
        .io_pins_qspi_dq_0_i_ival         (qspi_dq_ival[0]  ),
        .io_pins_qspi_dq_0_i_po           (/* UNCONNECTED */),
        .io_pins_qspi_dq_0_o_oval         (qspi_dq_oval[0]  ),
        .io_pins_qspi_dq_0_o_oe           (qspi_dq_oe[0]    ),
        .io_pins_qspi_dq_0_o_ie           (/* UNCONNECTED */),
        .io_pins_qspi_dq_1_i_ival         (qspi_dq_ival[1]  ),
        .io_pins_qspi_dq_1_i_po           (/* UNCONNECTED */),
        .io_pins_qspi_dq_1_o_oval         (qspi_dq_oval[1]  ),
        .io_pins_qspi_dq_1_o_oe           (qspi_dq_oe[1]    ),
        .io_pins_qspi_dq_1_o_ie           (/* UNCONNECTED */),
        .io_pins_qspi_dq_2_i_ival         (qspi_dq_ival[2]  ),
        .io_pins_qspi_dq_2_i_po           (/* UNCONNECTED */),
        .io_pins_qspi_dq_2_o_oval         (qspi_dq_oval[2]  ),
        .io_pins_qspi_dq_2_o_oe           (qspi_dq_oe[2]    ),
        .io_pins_qspi_dq_2_o_ie           (/* UNCONNECTED */),
        .io_pins_qspi_dq_3_i_ival         (qspi_dq_ival[3]  ),
        .io_pins_qspi_dq_3_i_po           (/* UNCONNECTED */),
        .io_pins_qspi_dq_3_o_oval         (qspi_dq_oval[3]  ),
        .io_pins_qspi_dq_3_o_oe           (qspi_dq_oe[3]    ),
        .io_pins_qspi_dq_3_o_ie           (/* UNCONNECTED */),
        .io_ndreset                       (/* UNCONNECTED */)
    );

endmodule